#define ILD_ROP 0x0040
#define   BP_PUSHBUTTON 1
#define   BP_RADIOBUTTON 2
#define   BP_CHECKBOX 3
#define   BP_GROUPBOX 4
#define   BP_USERBUTTON 5
#define   PBS_NORMAL 1
#define   PBS_HOT 2
#define   PBS_PRESSED 3
#define   PBS_DISABLED 4
#define   PBS_DEFAULTED 5
#define	DTT_GRAYED 1
