// Delete Window.vh

