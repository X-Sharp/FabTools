// Delete Window.vh

STATIC DEFINE DELETEWND_DELETEPB := 100 
STATIC DEFINE DELETEWND_CANCELPB := 101 
STATIC DEFINE DELETEWND_FILESGRP := 102 
STATIC DEFINE DELETEWND_SELECTRADIO := 103 
STATIC DEFINE DELETEWND_ALLRADIO := 104 
