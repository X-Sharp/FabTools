#define IDM_EmptyShellMenu_File_Paste_from_Clipboard_ID 17234
#define IDM_EmptyShellMenu "EmptyShellMenu"
#define IDA_EmptyShellMenu "EmptyShellMenu"
#define IDM_EmptyShellMenu_File_ID 17232
#define IDM_EmptyShellMenu_File_Open_ID 32001
#define IDM_EmptyShellMenu_File_Print_Setup_ID 17236
#define IDM_EmptyShellMenu_File_Exit_ID 17238
#define IDM_EmptyShellMenu_Help_ID 17239
#define IDM_EmptyShellMenu_Help_Index_ID 17240
#define IDM_EmptyShellMenu_Help_Using_help_ID 17241
#define IDM_EmptyShellMenu_Help_About_ID 32031
#define IDM_ImgViewShellMenu "ImgViewShellMenu"
#define IDA_ImgViewShellMenu "ImgViewShellMenu"
#define IDM_ImgViewShellMenu_File_ID 17108
#define IDM_ImgViewShellMenu_File_Open_ID 32001
#define IDM_ImgViewShellMenu_File_Save_As__ID 17110
#define IDM_ImgViewShellMenu_File_Close_ID 17111
#define IDM_ImgViewShellMenu_File_Print_ID 17113
#define IDM_ImgViewShellMenu_File_Print_Setup_ID 17114
#define IDM_ImgViewShellMenu_File_Send__ID 17116
#define IDM_ImgViewShellMenu_File_Exit_ID 17118
#define IDM_ImgViewShellMenu_Window_ID 17146
#define IDM_ImgViewShellMenu_Window_Cascade_ID 17147
#define IDM_ImgViewShellMenu_Window_Tile_ID 17148
#define IDM_ImgViewShellMenu_Window_Close_All_ID 17149
#define IDM_ImgViewShellMenu_Help_ID 17150
#define IDM_ImgViewShellMenu_Help_Index_ID 17151
#define IDM_ImgViewShellMenu_Help_Context_Help_ID 17152
#define IDM_ImgViewShellMenu_Help_Using_Help_ID 17153
#define IDM_ImgViewShellMenu_Help_About_ID 32031
#define IDM_ImgViewShellMenu_Image_ID 17122
#define IDM_ImgViewShellMenu_Image_Copy_ID 17123
#define IDM_ImgViewShellMenu_Image_Resize_ID 17128
#define IDM_ImgViewShellMenu_Image_Resize_Bilinear_ID 17129
#define IDM_ImgViewShellMenu_Image_Resize_Box_ID 17130
#define IDM_ImgViewShellMenu_Image_Resize_Gaussian_ID 17131
#define IDM_ImgViewShellMenu_Image_Resize_Hamming_ID 17132
#define IDM_ImgViewShellMenu_Image_Crop_ID 17133
#define IDM_ImgViewShellMenu_Image_Grayscale_ID 17134
#define IDM_ImgViewShellMenu_Image_Rotate_ID 17135
#define IDM_ImgViewShellMenu_Image_Invert_ID 17136
#define IDM_ImgViewShellMenu_Edit_ID 17119
#define IDM_ImgViewShellMenu_Edit_Copy_ID 17120
#define IDM_ImgViewShellMenu_Edit_Paste_ID 17121
#define IDM_ImgViewShellMenu_Image_Copy_No_Change_ID 17124
#define IDM_ImgViewShellMenu_Image_Copy__1_bpp_ID 17125
#define IDM_ImgViewShellMenu_Image_Copy__8_bpp_ID 17126
#define IDM_ImgViewShellMenu_Image_Copy__32_bpp_ID 17127
#define IDM_ImgViewShellMenu_Image_Contrast_ID 17141
#define IDM_ImgViewShellMenu_Image_Lightness_ID 17142
#define IDM_ImgViewShellMenu_Image_Intensity_ID 17143
#define IDM_ImgViewShellMenu_Image_EXIF_Data_ID 17145
#define IDM_ImgViewShellMenu_Image_Zoom_b2_ID 17138
#define IDM_ImgViewShellMenu_Image_Zoom__ID 17139
#define USE_CAPAINT .T. 
#define IDI_STANDARDICON 101
#define IDS_ERROR 65520
#define IDS_EXCHANGE_NOT_INSTALLED 65521
#define IDS_SAVE 65522
