// Wnd ImgView.vh

#define HELPABOUT_PUSHBUTTON1 (104 )
#define MAILDLG_RICHEDIT1 (100 )
#define MAILDLG_PBSEND (102 )
#define MAILDLG_PBCANCEL (101 )
#define HELPABOUT_FIXEDICON1 (100 )
#define HELPABOUT_FIXEDTEXT1 (101 )
#define HELPABOUT_FIXEDTEXT2 (102 )
#define HELPABOUT_FIXEDTEXT3 (103 )
#define PROGRESS_PROGRESSBAR1 (100 )
#define INPUTBOX_VALUE1TXT (100 )
#define INPUTBOX_VALUE1 (101 )
#define INPUTBOX_VALUE2 (102 )
#define INPUTBOX_VALUE2TXT (103 )
#define INPUTBOX_VALUE3TXT (104 )
#define INPUTBOX_VALUE3 (105 )
#define INPUTBOX_VALUE4 (106 )
#define INPUTBOX_VALUE4TXT (107 )
#define INPUTBOX_OKPB (108 )
#define INPUTBOX_CANCELPB (109 )
