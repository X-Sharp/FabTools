// Dlg EXIF.vh

#define EXIFDLG_CLOSEPB (100 )
#define EXIFDLG_EXIFLISTVIEW (101 )
