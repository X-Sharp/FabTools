// Dlg Progress.vh

#define PROGRESS_PROGRESSBAR1 (100 )
