// Extract Window.vh

#define SELECTPATH_OKPB (100 )
#define SELECTPATH_CANCELPB (101 )
