// Dlg EXIF.vh

