// Dlg About.vh

#define HELPABOUT_FIXEDICON1 (100 )
#define HELPABOUT_FIXEDTEXT1 (101 )
#define HELPABOUT_FIXEDTEXT2 (102 )
#define HELPABOUT_PUSHBUTTON1 (103 )
