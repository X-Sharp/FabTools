#define IDM_ListMenu "ListMenu"
#define IDA_ListMenu "ListMenu"
#define IDM_ListMenu_Dummy_ID 18325
#define IDM_ListMenu_Dummy_Select_All_ID 18326
#define IDM_ListMenu_Dummy_Deselect_All_ID 18327
#define IDM_ListMenu_Dummy_Add_ID 18329
#define IDM_ListMenu_Dummy_Extract_ID 18330
#define IDM_ListMenu_Dummy_Delete_ID 18331
#define IDM_StandardShellMenu "StandardShellMenu"
#define IDA_StandardShellMenu "StandardShellMenu"
#define IDM_StandardShellMenu_File_ID 15097
#define IDM_StandardShellMenu_File_Open_ID 32001
#define IDM_StandardShellMenu_File_Close_ID 15099
#define IDM_StandardShellMenu_File_Print_Setup_ID 15102
#define IDM_StandardShellMenu_File_Send__ID 15104
#define IDM_StandardShellMenu_File_Exit_ID 15106
#define IDM_StandardShellMenu_Edit_ID 15107
#define IDM_StandardShellMenu_Edit_Cut_ID 15108
#define IDM_StandardShellMenu_Edit_Copy_ID 15109
#define IDM_StandardShellMenu_Edit_Paste_ID 15110
#define IDM_StandardShellMenu_Edit_Insert_Record_ID 15112
#define IDM_StandardShellMenu_Edit_Delete_Record_ID 15113
#define IDM_StandardShellMenu_Edit_Go_To_Top_ID 15115
#define IDM_StandardShellMenu_Edit_Previous_ID 15116
#define IDM_StandardShellMenu_Edit_Next_ID 15117
#define IDM_StandardShellMenu_Edit_Go_To_Bottom_ID 15118
#define IDM_StandardShellMenu_View_ID 15119
#define IDM_StandardShellMenu_View_Form_ID 15120
#define IDM_StandardShellMenu_View_Table_ID 15121
#define IDM_StandardShellMenu_Window_ID 15122
#define IDM_StandardShellMenu_Window_Cascade_ID 15123
#define IDM_StandardShellMenu_Window_Tile_ID 15124
#define IDM_StandardShellMenu_Window_Close_All_ID 15125
#define IDM_StandardShellMenu_Help_ID 15126
#define IDM_StandardShellMenu_Help_Index_ID 15127
#define IDM_StandardShellMenu_Help_Context_Help_ID 15128
#define IDM_StandardShellMenu_Help_Using_Help_ID 15129
#define IDM_StandardShellMenu_Help_About_ID 32031
#define IDM_StandardShellMenu_File_Print_ID 15101
#define IDM_MenuStd "MenuStd"
#define IDA_MenuStd "MenuStd"
#define IDM_MenuStd_FabZip_ID 15337
#define IDM_MenuStd_FabZip_Test_ID 32001
#define IDM_MenuStd_FabZip_Exit_ID 15340
#define IDM_MenuStd_Help_ID 15341
#define IDM_MenuStd_Help_About_ID 32031
