// Add Window.vh

STATIC DEFINE ADDWND_FIXEDTEXT1 := 117 
STATIC DEFINE ADDWND_DOITPB := 114 
STATIC DEFINE ADDWND_CANCELPB := 116 
STATIC DEFINE ADDWND_SELECTPB := 101 
STATIC DEFINE ADDWND_FIXEDTEXT2 := 118 
STATIC DEFINE ADDWND_ACTIONCOMBO := 102 
STATIC DEFINE ADDWND_FIXEDTEXT3 := 119 
STATIC DEFINE ADDWND_LEVELSLIDER := 103 
STATIC DEFINE ADDWND_FIXEDTEXT4 := 120 
STATIC DEFINE ADDWND_FIXEDTEXT5 := 121 
STATIC DEFINE ADDWND_FILES := 100 
STATIC DEFINE ADDWND_WILDCARDSPB := 115 
STATIC DEFINE ADDWND_FOLDERSGRP := 122 
STATIC DEFINE ADDWND_RECURSECHK := 106 
STATIC DEFINE ADDWND_DIRINFOCHK := 107 
STATIC DEFINE ADDWND_SYSTEMCHK := 105 
STATIC DEFINE ADDWND_DOSFORMATCHK := 104 
STATIC DEFINE ADDWND_FORMATCHK := 110 
STATIC DEFINE ADDWND_FIXEDTEXT6 := 123 
STATIC DEFINE ADDWND_MINFREESIZE := 113 
STATIC DEFINE ADDWND_DISKSIZEGRP := 124 
STATIC DEFINE ADDWND_FIXEDTEXT7 := 125 
STATIC DEFINE ADDWND_MINDISK1 := 112 
STATIC DEFINE ADDWND_FIXEDTEXT8 := 126 
STATIC DEFINE ADDWND_MAXSIZE := 111 
STATIC DEFINE ADDWND_DISKSPANNINGGRP := 108 
STATIC DEFINE ADDWND_SPANNINGCHK := 109 
