#define GRADIENT_FILL_RECT_H 0
#define GRADIENT_FILL_RECT_V 1
#define GRADIENT_FILL_RECT_TRIANGLE 2
