// Dlg About.vh

