// Test Window.vh

STATIC DEFINE FABZIPTEST1_OKPB := 109 
STATIC DEFINE FABZIPTEST1_ZIP_CONTROL := 110 
STATIC DEFINE FABZIPTEST1_ZIPFILENAME := 100 
STATIC DEFINE FABZIPTEST1_ZIPLIST := 111 
STATIC DEFINE FABZIPTEST1_GROUPBOX1 := 114 
STATIC DEFINE FABZIPTEST1_EXTRACTPB := 105 
STATIC DEFINE FABZIPTEST1_FPROCESS := 116 
STATIC DEFINE FABZIPTEST1_DLLMSG := 112 
STATIC DEFINE FABZIPTEST1_ADDPB := 104 
STATIC DEFINE FABZIPTEST1_DELETEPB := 106 
STATIC DEFINE FABZIPTEST1_CANCELPB := 117 
STATIC DEFINE FABZIPTEST1_PROCESSGRP := 118 
STATIC DEFINE FABZIPTEST1_OPENPB := 101 
STATIC DEFINE FABZIPTEST1_CREATEPB := 102 
STATIC DEFINE FABZIPTEST1_PASSCHK := 103 
STATIC DEFINE FABZIPTEST1_CONVERTPB := 107 
STATIC DEFINE FABZIPTEST1_EXTRACTBAR := 115 
STATIC DEFINE FABZIPTEST1_COMMENTPB := 108 
STATIC DEFINE FABZIPTEST1_TOTALFILESBAR := 120 
STATIC DEFINE FABZIPTEST1_TOTALSIZEBAR := 119 
STATIC DEFINE FABZIPTEST1_FABZIPMSG := 113 
STATIC DEFINE FABZIPTEST1_ZIPMESSAGES := 121 
