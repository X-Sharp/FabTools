// Add Window.vh

