Define IDM_ListMenu := "ListMenu"
Define IDA_ListMenu := "ListMenu"
Define IDM_ListMenu_Dummy_ID := 18325
Define IDM_ListMenu_Dummy_Select_All_ID := 18326
Define IDM_ListMenu_Dummy_Deselect_All_ID := 18327
Define IDM_ListMenu_Dummy_Add_ID := 18329
Define IDM_ListMenu_Dummy_Extract_ID := 18330
Define IDM_ListMenu_Dummy_Delete_ID := 18331
Define IDM_StandardShellMenu := "StandardShellMenu"
Define IDA_StandardShellMenu := "StandardShellMenu"
Define IDM_StandardShellMenu_File_ID := 15097
Define IDM_StandardShellMenu_File_Open_ID := 32001
Define IDM_StandardShellMenu_File_Close_ID := 15099
Define IDM_StandardShellMenu_File_Print_Setup_ID := 15102
Define IDM_StandardShellMenu_File_Send__ID := 15104
Define IDM_StandardShellMenu_File_Exit_ID := 15106
Define IDM_StandardShellMenu_Edit_ID := 15107
Define IDM_StandardShellMenu_Edit_Cut_ID := 15108
Define IDM_StandardShellMenu_Edit_Copy_ID := 15109
Define IDM_StandardShellMenu_Edit_Paste_ID := 15110
Define IDM_StandardShellMenu_Edit_Insert_Record_ID := 15112
Define IDM_StandardShellMenu_Edit_Delete_Record_ID := 15113
Define IDM_StandardShellMenu_Edit_Go_To_Top_ID := 15115
Define IDM_StandardShellMenu_Edit_Previous_ID := 15116
Define IDM_StandardShellMenu_Edit_Next_ID := 15117
Define IDM_StandardShellMenu_Edit_Go_To_Bottom_ID := 15118
Define IDM_StandardShellMenu_View_ID := 15119
Define IDM_StandardShellMenu_View_Form_ID := 15120
Define IDM_StandardShellMenu_View_Table_ID := 15121
Define IDM_StandardShellMenu_Window_ID := 15122
Define IDM_StandardShellMenu_Window_Cascade_ID := 15123
Define IDM_StandardShellMenu_Window_Tile_ID := 15124
Define IDM_StandardShellMenu_Window_Close_All_ID := 15125
Define IDM_StandardShellMenu_Help_ID := 15126
Define IDM_StandardShellMenu_Help_Index_ID := 15127
Define IDM_StandardShellMenu_Help_Context_Help_ID := 15128
Define IDM_StandardShellMenu_Help_Using_Help_ID := 15129
Define IDM_StandardShellMenu_Help_About_ID := 32031
Define IDM_StandardShellMenu_File_Print_ID := 15101
Define IDM_MenuStd := "MenuStd"
Define IDA_MenuStd := "MenuStd"
Define IDM_MenuStd_FabZip_ID := 15337
Define IDM_MenuStd_FabZip_Test_ID := 32001
Define IDM_MenuStd_FabZip_Exit_ID := 15340
Define IDM_MenuStd_Help_ID := 15341
Define IDM_MenuStd_Help_About_ID := 32031
