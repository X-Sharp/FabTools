// Test Window.vh

