// Dlg Progress.vh

