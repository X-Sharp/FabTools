// Dlg Input.vh

