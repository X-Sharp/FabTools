// About.vh

STATIC DEFINE HELPABOUT_FIXEDICON1 := 102 
STATIC DEFINE HELPABOUT_FIXEDTEXT2 := 101 
STATIC DEFINE HELPABOUT_FIXEDTEXT3 := 104 
STATIC DEFINE HELPABOUT_OKPB := 105 
STATIC DEFINE HELPABOUT_DLLINFOPB := 100 
STATIC DEFINE HELPABOUT_FABZIPVERSION := 103 
