#define TIFF_DEFAULT 0
#define TIFF_CMYK (0x0001 )
#define TIFF_PACKBITS (0x0100 )
#define TIFF_DEFLATE (0x0200 )
#define TIFF_ADOBE_DEFLATE (0x0400 )
#define TIFF_NONE (0x0800 )
#define TIFF_CCITTFAX3 (0x1000 )
#define TIFF_CCITTFAX4 (0x2000 )
#define TIFF_LZW (0x4000 )
#define TIFF_JPEG (0x8000 )
#define	    COMPRESSION_PACKBITS (0x0100 )
#define	    COMPRESSION_NONE (0x0800 )
#define	    COMPRESSION_CCITTFAX3 (0x1000 )
#define	    COMPRESSION_CCITTFAX4 (0x2000 )
#define	    COMPRESSION_LZW (0x4000 )
#define	    COMPRESSION_JPEG (0x8000 )
#define	    COMPRESSION_DEFLATE (0x0200 )
#define     COMPRESSION_ADOBE_DEFLATE (0x0400 )
#define EXIF_MODEL_COMMENTS 0
#define EXIF_MODEL_MAIN FREE_IMAGE_MDMODEL.FIMD_EXIF_MAIN
#define EXIF_MODEL_EXIF FREE_IMAGE_MDMODEL.FIMD_EXIF_EXIF
#define EXIF_MODEL_GPS FREE_IMAGE_MDMODEL.FIMD_EXIF_GPS
#define EXIF_MODEL_MAKERNOTE FREE_IMAGE_MDMODEL.FIMD_EXIF_MAKERNOTE
#define EXIF_MODEL_INTEROP 5
#define EXIF_MODEL_IPTC 6
#define EXIF_MODEL_XMP 7
#define EXIF_MODEL_GEOTIFF 8
#define EXIF_MODEL_ANIMATION 9
#define EXIF_MODEL_CUSTOM 10
#define EXIF_MODEL_NONE (-1)
