// Extract Window.vh

STATIC DEFINE SELECTPATH_OKPB := 100 
STATIC DEFINE SELECTPATH_CANCELPB := 101 
STATIC DEFINE EXTRACTWND_SELECTRADIO := 103 
STATIC DEFINE EXTRACTWND_ALLRADIO := 104 
STATIC DEFINE EXTRACTWND_FILESGROUP := 102 
STATIC DEFINE EXTRACTWND_DIRNAME := 110 
STATIC DEFINE EXTRACTWND_OVERWRITE := 109 
STATIC DEFINE EXTRACTWND_SLEDIR := 100 
STATIC DEFINE EXTRACTWND_PBOK := 111 
STATIC DEFINE EXTRACTWND_PBCANCEL := 112 
STATIC DEFINE EXTRACTWND_FOLDERSTV := 101 
STATIC DEFINE EXTRACTWND_NORMALBTN := 106 
STATIC DEFINE EXTRACTWND_FRESHENBTN := 107 
STATIC DEFINE EXTRACTWND_UPDATEBTN := 108 
STATIC DEFINE EXTRACTWND_EXTRACTGROUP := 105 
STATIC DEFINE EXTRACTWND_FIXEDTEXT1 := 113 
STATIC DEFINE EXTRACTWND_FIXEDTEXT2 := 114 
