// SFX Window.vh

STATIC DEFINE SFXWND_OKPB := 100 
STATIC DEFINE SFXWND_HELPPB := 101 
STATIC DEFINE SFXWND_SFXCAPTION := 102 
STATIC DEFINE SFXWND_FIXEDTEXT1 := 103 
STATIC DEFINE SFXWND_FIXEDTEXT2 := 105 
STATIC DEFINE SFXWND_FIXEDTEXT3 := 107 
STATIC DEFINE SFXWND_CMDCHK := 108 
STATIC DEFINE SFXWND_FILESCHK := 109 
STATIC DEFINE SFXWND_FIXEDTEXT4 := 110 
STATIC DEFINE SFXWND_OVERCHK := 111 
STATIC DEFINE SFXWND_SFXDEFAULTDIR := 104 
STATIC DEFINE SFXWND_SFXCOMMANDLINE := 106 
STATIC DEFINE SFXWND_OVERCOMBO := 112 
STATIC DEFINE SFXWND_CANCELPB := 113 
