// SFX Window.vh

